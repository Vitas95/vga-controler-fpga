module font_memory (
  input clock,
  input reset
);



endmodule